-- Created by Eduardo Flores in fulfillment of his Bachellor's degree Thesis.


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.ldpc_encoder_pac.ALL;

ENTITY addresses IS
  PORT( slot                              :   IN    std_logic_vector(7 DOWNTO 0);  -- uint8
        counter                           :   IN    std_logic_vector(8 DOWNTO 0);  -- ufix9
        q_factor                          :   IN    std_logic_vector(7 DOWNTO 0);  -- uint8
        addresses_1                       :   OUT   vector_of_std_logic_vector16(0 TO 11)  -- uint16 [12]
        );
END addresses;


ARCHITECTURE rtl OF addresses IS

  -- Constants
  CONSTANT nc                             : matrix_of_signed16(0 TO 134, 0 TO 11) := 
    (( to_signed(16#0000#, 16), to_signed(16#18F1#, 16), to_signed(16#1EDD#, 16), to_signed(16#3913#, 16),
     to_signed(16#344D#, 16), to_signed(16#2BC0#, 16), to_signed(16#0CB4#, 16), to_signed(16#147B#, 16),
     to_signed(16#09C8#, 16), to_signed(16#0AA2#, 16), to_signed(16#0335#, 16), to_signed(16#1CCE#, 16) ),
     ( to_signed(16#0001#, 16), to_signed(16#2C5F#, 16), to_signed(16#0A8A#, 16), to_signed(16#0165#, 16),
     to_signed(16#3600#, 16), to_signed(16#31E4#, 16), to_signed(16#1C4C#, 16), to_signed(16#1A60#, 16),
     to_signed(16#3BCE#, 16), to_signed(16#0354#, 16), to_signed(16#07D1#, 16), to_signed(16#2C99#, 16) ),
     ( to_signed(16#0002#, 16), to_signed(16#1EB6#, 16), to_signed(16#1F29#, 16), to_signed(16#18B1#, 16),
     to_signed(16#352C#, 16), to_signed(16#2FA5#, 16), to_signed(16#3871#, 16), to_signed(16#3B21#, 16),
     to_signed(16#3624#, 16), to_signed(16#06AC#, 16), to_signed(16#18FF#, 16), to_signed(16#3484#, 16) ),
     ( to_signed(16#0003#, 16), to_signed(16#0618#, 16), to_signed(16#2E1C#, 16), to_signed(16#1B3F#, 16),
     to_signed(16#33EC#, 16), to_signed(16#0E3E#, 16), to_signed(16#0EE4#, 16), to_signed(16#2244#, 16),
     to_signed(16#1C8A#, 16), to_signed(16#16A3#, 16), to_signed(16#37F7#, 16), to_signed(16#1EBA#, 16) ),
     ( to_signed(16#0004#, 16), to_signed(16#1DCA#, 16), to_signed(16#2C8F#, 16), to_signed(16#3907#, 16),
     to_signed(16#25D9#, 16), to_signed(16#065C#, 16), to_signed(16#0841#, 16), to_signed(16#2A39#, 16),
     to_signed(16#2443#, 16), to_signed(16#04CE#, 16), to_signed(16#3B89#, 16), to_signed(16#1306#, 16) ),
     ( to_signed(16#0005#, 16), to_signed(16#064A#, 16), to_signed(16#1643#, 16), to_signed(16#3E04#, 16),
     to_signed(16#24E6#, 16), to_signed(16#30E3#, 16), to_signed(16#0578#, 16), to_signed(16#189F#, 16),
     to_signed(16#1523#, 16), to_signed(16#3765#, 16), to_signed(16#3665#, 16), to_signed(16#1CBE#, 16) ),
     ( to_signed(16#0006#, 16), to_signed(16#0FDB#, 16), to_signed(16#2284#, 16), to_signed(16#0D4D#, 16),
     to_signed(16#1EAD#, 16), to_signed(16#1F38#, 16), to_signed(16#3BE8#, 16), to_signed(16#1752#, 16),
     to_signed(16#2880#, 16), to_signed(16#2826#, 16), to_signed(16#25CB#, 16), to_signed(16#122B#, 16) ),
     ( to_signed(16#0007#, 16), to_signed(16#1159#, 16), to_signed(16#0F7B#, 16), to_signed(16#23C1#, 16),
     to_signed(16#083D#, 16), to_signed(16#318B#, 16), to_signed(16#1D23#, 16), to_signed(16#2EFE#, 16),
     to_signed(16#2FBD#, 16), to_signed(16#0275#, 16), to_signed(16#3B6C#, 16), to_signed(16#0196#, 16) ),
     ( to_signed(16#0008#, 16), to_signed(16#1777#, 16), to_signed(16#20DB#, 16), to_signed(16#168B#, 16),
     to_signed(16#0DA9#, 16), to_signed(16#021F#, 16), to_signed(16#377A#, 16), to_signed(16#036B#, 16),
     to_signed(16#23E2#, 16), to_signed(16#185B#, 16), to_signed(16#3654#, 16), to_signed(16#0DEB#, 16) ),
     ( to_signed(16#0009#, 16), to_signed(16#0CA0#, 16), to_signed(16#19E1#, 16), to_signed(16#12BB#, 16),
     to_signed(16#0222#, 16), to_signed(16#2635#, 16), to_signed(16#0817#, 16), to_signed(16#1C90#, 16),
     to_signed(16#0D47#, 16), to_signed(16#1C52#, 16), to_signed(16#1344#, 16), to_signed(16#316C#, 16) ),
     ( to_signed(16#000A#, 16), to_signed(16#2274#, 16), to_signed(16#2768#, 16), to_signed(16#2B52#, 16),
     to_signed(16#1B9D#, 16), to_signed(16#19B9#, 16), to_signed(16#334E#, 16), to_signed(16#27AE#, 16),
     to_signed(16#1C0F#, 16), to_signed(16#01E8#, 16), to_signed(16#1D1F#, 16), to_signed(16#2416#, 16) ),
     ( to_signed(16#000B#, 16), to_signed(16#076F#, 16), to_signed(16#2A42#, 16), to_signed(16#0077#, 16),
     to_signed(16#00D7#, 16), to_signed(16#1D86#, 16), to_signed(16#2B26#, 16), to_signed(16#2977#, 16),
     to_signed(16#2D19#, 16), to_signed(16#39C0#, 16), to_signed(16#1F19#, 16), to_signed(16#3D03#, 16) ),
     ( to_signed(16#000C#, 16), to_signed(16#0E47#, 16), to_signed(16#2220#, 16), to_signed(16#1335#, 16),
     to_signed(16#3E02#, 16), to_signed(16#1409#, 16), to_signed(16#0856#, 16), to_signed(16#3E48#, 16),
     to_signed(16#39B0#, 16), to_signed(16#1BEE#, 16), to_signed(16#0A84#, 16), to_signed(16#05BD#, 16) ),
     ( to_signed(16#000D#, 16), to_signed(16#207C#, 16), to_signed(16#0EEC#, 16), to_signed(16#01F9#, 16),
     to_signed(16#22DB#, 16), to_signed(16#1A65#, 16), to_signed(16#0326#, 16), to_signed(16#1F15#, 16),
     to_signed(16#1078#, 16), to_signed(16#3CE5#, 16), to_signed(16#33BC#, 16), to_signed(16#0A3E#, 16) ),
     ( to_signed(16#000E#, 16), to_signed(16#387F#, 16), to_signed(16#12F4#, 16), to_signed(16#3D75#, 16),
     to_signed(16#0BE1#, 16), to_signed(16#2BB9#, 16), to_signed(16#323C#, 16), to_signed(16#3569#, 16),
     to_signed(16#1FD8#, 16), to_signed(16#1997#, 16), to_signed(16#3B04#, 16), to_signed(16#2236#, 16) ),
     ( to_signed(16#000F#, 16), to_signed(16#0C4D#, 16), to_signed(16#2ECD#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0010#, 16), to_signed(16#3468#, 16), to_signed(16#1AFA#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0011#, 16), to_signed(16#332A#, 16), to_signed(16#3428#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0012#, 16), to_signed(16#07D9#, 16), to_signed(16#387C#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0013#, 16), to_signed(16#1C27#, 16), to_signed(16#10DA#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0014#, 16), to_signed(16#0CF0#, 16), to_signed(16#0F69#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0015#, 16), to_signed(16#1142#, 16), to_signed(16#1868#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0016#, 16), to_signed(16#0A6D#, 16), to_signed(16#3697#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0017#, 16), to_signed(16#1D93#, 16), to_signed(16#233F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0018#, 16), to_signed(16#375C#, 16), to_signed(16#0B97#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0019#, 16), to_signed(16#1C67#, 16), to_signed(16#1BE2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001A#, 16), to_signed(16#17F7#, 16), to_signed(16#3566#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001B#, 16), to_signed(16#1D42#, 16), to_signed(16#38DF#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001C#, 16), to_signed(16#21D1#, 16), to_signed(16#09A2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001D#, 16), to_signed(16#2197#, 16), to_signed(16#3222#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001E#, 16), to_signed(16#0D8E#, 16), to_signed(16#0C50#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001F#, 16), to_signed(16#365D#, 16), to_signed(16#110D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0020#, 16), to_signed(16#1788#, 16), to_signed(16#35A2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0021#, 16), to_signed(16#2ADD#, 16), to_signed(16#3766#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0022#, 16), to_signed(16#09A0#, 16), to_signed(16#336F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0023#, 16), to_signed(16#14A1#, 16), to_signed(16#3AC9#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0024#, 16), to_signed(16#044F#, 16), to_signed(16#0739#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0025#, 16), to_signed(16#080A#, 16), to_signed(16#042D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0026#, 16), to_signed(16#25B6#, 16), to_signed(16#17CF#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0027#, 16), to_signed(16#37E7#, 16), to_signed(16#1DF3#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0028#, 16), to_signed(16#3D01#, 16), to_signed(16#1FD2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0029#, 16), to_signed(16#11EC#, 16), to_signed(16#2BD2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002A#, 16), to_signed(16#355C#, 16), to_signed(16#1863#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002B#, 16), to_signed(16#2182#, 16), to_signed(16#1EC2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002C#, 16), to_signed(16#2DDD#, 16), to_signed(16#0A7E#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0000#, 16), to_signed(16#03FE#, 16), to_signed(16#04F0#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0001#, 16), to_signed(16#313C#, 16), to_signed(16#26ED#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0002#, 16), to_signed(16#2019#, 16), to_signed(16#0A93#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0003#, 16), to_signed(16#0C54#, 16), to_signed(16#2E11#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0004#, 16), to_signed(16#0162#, 16), to_signed(16#05EA#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0005#, 16), to_signed(16#1B42#, 16), to_signed(16#36EA#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0006#, 16), to_signed(16#1EF2#, 16), to_signed(16#3ECF#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0007#, 16), to_signed(16#3AEF#, 16), to_signed(16#2F6A#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0008#, 16), to_signed(16#13BD#, 16), to_signed(16#1946#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0009#, 16), to_signed(16#318F#, 16), to_signed(16#3A54#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000A#, 16), to_signed(16#3C62#, 16), to_signed(16#06E3#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000B#, 16), to_signed(16#1FB9#, 16), to_signed(16#06B9#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000C#, 16), to_signed(16#308F#, 16), to_signed(16#0225#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000D#, 16), to_signed(16#1021#, 16), to_signed(16#1BB3#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000E#, 16), to_signed(16#0592#, 16), to_signed(16#20DF#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000F#, 16), to_signed(16#2637#, 16), to_signed(16#1DB4#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0010#, 16), to_signed(16#1897#, 16), to_signed(16#2C41#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0011#, 16), to_signed(16#0581#, 16), to_signed(16#2F1D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0012#, 16), to_signed(16#1F81#, 16), to_signed(16#237F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0013#, 16), to_signed(16#0B66#, 16), to_signed(16#20F6#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0014#, 16), to_signed(16#050D#, 16), to_signed(16#3723#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0015#, 16), to_signed(16#0F52#, 16), to_signed(16#361B#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0016#, 16), to_signed(16#0F0B#, 16), to_signed(16#0FA0#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0017#, 16), to_signed(16#16E9#, 16), to_signed(16#06E8#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0018#, 16), to_signed(16#0A5F#, 16), to_signed(16#3A6D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0019#, 16), to_signed(16#15BD#, 16), to_signed(16#18BC#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001A#, 16), to_signed(16#10CF#, 16), to_signed(16#3157#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001B#, 16), to_signed(16#2D85#, 16), to_signed(16#2FCC#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001C#, 16), to_signed(16#3E99#, 16), to_signed(16#1DD0#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001D#, 16), to_signed(16#122F#, 16), to_signed(16#3730#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001E#, 16), to_signed(16#2570#, 16), to_signed(16#3343#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001F#, 16), to_signed(16#36A3#, 16), to_signed(16#257D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0020#, 16), to_signed(16#3C31#, 16), to_signed(16#2F4E#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0021#, 16), to_signed(16#2232#, 16), to_signed(16#3C82#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0022#, 16), to_signed(16#1CF8#, 16), to_signed(16#3BDD#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0023#, 16), to_signed(16#0B5D#, 16), to_signed(16#3CBD#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0024#, 16), to_signed(16#0BB3#, 16), to_signed(16#2041#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0025#, 16), to_signed(16#24BE#, 16), to_signed(16#12B7#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0026#, 16), to_signed(16#2B67#, 16), to_signed(16#12F6#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0027#, 16), to_signed(16#0AFC#, 16), to_signed(16#2149#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0028#, 16), to_signed(16#211C#, 16), to_signed(16#397D#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0029#, 16), to_signed(16#1E8C#, 16), to_signed(16#3C00#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002A#, 16), to_signed(16#049B#, 16), to_signed(16#1F03#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002B#, 16), to_signed(16#0935#, 16), to_signed(16#21E6#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002C#, 16), to_signed(16#1E17#, 16), to_signed(16#1848#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0000#, 16), to_signed(16#0D95#, 16), to_signed(16#1B9B#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0001#, 16), to_signed(16#0F5B#, 16), to_signed(16#3615#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0002#, 16), to_signed(16#1DFB#, 16), to_signed(16#3263#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0003#, 16), to_signed(16#06DA#, 16), to_signed(16#1FFB#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0004#, 16), to_signed(16#1E69#, 16), to_signed(16#0578#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0005#, 16), to_signed(16#23FD#, 16), to_signed(16#1703#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0006#, 16), to_signed(16#09BE#, 16), to_signed(16#1E17#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0007#, 16), to_signed(16#0A10#, 16), to_signed(16#1EDE#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0008#, 16), to_signed(16#12D5#, 16), to_signed(16#3D42#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0009#, 16), to_signed(16#28BA#, 16), to_signed(16#2E9F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000A#, 16), to_signed(16#0712#, 16), to_signed(16#0388#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000B#, 16), to_signed(16#2C44#, 16), to_signed(16#2430#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000C#, 16), to_signed(16#2C30#, 16), to_signed(16#0DF2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000D#, 16), to_signed(16#3A44#, 16), to_signed(16#0A5A#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000E#, 16), to_signed(16#1DFF#, 16), to_signed(16#1EA2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#000F#, 16), to_signed(16#17C9#, 16), to_signed(16#331C#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0010#, 16), to_signed(16#0F62#, 16), to_signed(16#0ABF#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0011#, 16), to_signed(16#213D#, 16), to_signed(16#1228#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0012#, 16), to_signed(16#2FAC#, 16), to_signed(16#22D5#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0013#, 16), to_signed(16#1675#, 16), to_signed(16#309B#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0014#, 16), to_signed(16#3145#, 16), to_signed(16#114F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0015#, 16), to_signed(16#0540#, 16), to_signed(16#0FAE#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0016#, 16), to_signed(16#2128#, 16), to_signed(16#361A#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0017#, 16), to_signed(16#06C2#, 16), to_signed(16#3A30#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0018#, 16), to_signed(16#3A5E#, 16), to_signed(16#1BD6#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0019#, 16), to_signed(16#3A87#, 16), to_signed(16#229F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001A#, 16), to_signed(16#19B2#, 16), to_signed(16#2174#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001B#, 16), to_signed(16#1353#, 16), to_signed(16#018C#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001C#, 16), to_signed(16#0129#, 16), to_signed(16#3205#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001D#, 16), to_signed(16#3636#, 16), to_signed(16#1A24#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001E#, 16), to_signed(16#2E51#, 16), to_signed(16#2BB2#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#001F#, 16), to_signed(16#383B#, 16), to_signed(16#2CE5#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0020#, 16), to_signed(16#3F11#, 16), to_signed(16#2FDB#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0021#, 16), to_signed(16#3496#, 16), to_signed(16#1D04#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0022#, 16), to_signed(16#38BE#, 16), to_signed(16#333F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0023#, 16), to_signed(16#09E7#, 16), to_signed(16#2BEB#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0024#, 16), to_signed(16#1941#, 16), to_signed(16#3192#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0025#, 16), to_signed(16#1AD8#, 16), to_signed(16#2476#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0026#, 16), to_signed(16#3C0B#, 16), to_signed(16#36C7#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0027#, 16), to_signed(16#1FA5#, 16), to_signed(16#27CB#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0028#, 16), to_signed(16#2EBB#, 16), to_signed(16#12F0#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#0029#, 16), to_signed(16#3B15#, 16), to_signed(16#17E7#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002A#, 16), to_signed(16#1F73#, 16), to_signed(16#3881#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002B#, 16), to_signed(16#2B83#, 16), to_signed(16#142F#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ),
     ( to_signed(16#002C#, 16), to_signed(16#0B43#, 16), to_signed(16#38B9#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16),
     to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16), to_signed(16#3F48#, 16) ));  -- int16 [135x12]

  -- Signals
  SIGNAL slot_unsigned                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL counter_unsigned                 : unsigned(8 DOWNTO 0);  -- ufix9
  SIGNAL q_factor_unsigned                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL addresses_tmp                    : vector_of_unsigned16(0 TO 11);  -- uint16 [12]

BEGIN
  slot_unsigned <= unsigned(slot);

  counter_unsigned <= unsigned(counter);

  q_factor_unsigned <= unsigned(q_factor);

  addresses_2_output : PROCESS (counter_unsigned, q_factor_unsigned, slot_unsigned)
    VARIABLE buffer_rsvd : vector_of_unsigned16(0 TO 11);
    VARIABLE a : vector_of_unsigned16(0 TO 11);
    VARIABLE b : unsigned(7 DOWNTO 0);
    VARIABLE c : unsigned(16 DOWNTO 0);
    VARIABLE sub_cast : vector_of_signed32(0 TO 11);
    VARIABLE buffer_rsvd_0 : vector_of_unsigned16(0 TO 11);
  BEGIN
    --MATLAB Function 'ldpc_encoder/address_calculator/addresses'
    b := q_factor_unsigned;
    c := counter_unsigned * b;

    FOR t_0 IN 0 TO 11 LOOP
      sub_cast(t_0) := signed(resize(slot_unsigned, 32));
      a(t_0) := unsigned(nc(to_integer(sub_cast(t_0) - 1), t_0));
      buffer_rsvd(t_0) := resize(resize(a(t_0), 18) + resize(c, 18), 16);
      IF buffer_rsvd(t_0) >= to_unsigned(16#00003F48#, 16) THEN 
        buffer_rsvd_0(t_0) := to_unsigned(16#3F48#, 16);
      ELSE 
        buffer_rsvd_0(t_0) := to_unsigned(16#0000#, 16);
      END IF;
      addresses_tmp(t_0) <= buffer_rsvd(t_0) - buffer_rsvd_0(t_0);
    END LOOP;

  END PROCESS addresses_2_output;


  addresses_1(0) <= std_logic_vector(addresses_tmp(0));
  addresses_1(1) <= std_logic_vector(addresses_tmp(1));
  addresses_1(2) <= std_logic_vector(addresses_tmp(2));
  addresses_1(3) <= std_logic_vector(addresses_tmp(3));
  addresses_1(4) <= std_logic_vector(addresses_tmp(4));
  addresses_1(5) <= std_logic_vector(addresses_tmp(5));
  addresses_1(6) <= std_logic_vector(addresses_tmp(6));
  addresses_1(7) <= std_logic_vector(addresses_tmp(7));
  addresses_1(8) <= std_logic_vector(addresses_tmp(8));
  addresses_1(9) <= std_logic_vector(addresses_tmp(9));
  addresses_1(10) <= std_logic_vector(addresses_tmp(10));
  addresses_1(11) <= std_logic_vector(addresses_tmp(11));

END rtl;

